module number_rom
(
	input [7:0] address,
	output [7:0] data
);

	parameter[0:79][7:0] ROM = {
	
		8'b00000000, //
		8'b00011000, //   ██   
		8'b00100100, //  █  █  
		8'b01000010, // █    █ 
		8'b01000010, // █    █ 
		8'b00100100, //  █  █  
		8'b00011000, //   ██
		8'b00000000, //
		
		8'b00000000, // 
		8'b00001000, //     █  
		8'b00011000, //    ██   
		8'b00001000, //     █
		8'b00001000, //     █
		8'b00001000, //     █
		8'b00011100, //    ███
		8'b00000000, // 
		
		8'b00000000, // 
		8'b00011100, //    ███  
		8'b00100010, //   █   █ 
		8'b00000010, //       █
		8'b00011100, //    ███  
		8'b00100000, //   █     
		8'b00111110, //   █████ 
		8'b00000000, // 
		
		8'b00000000, //
		8'b00111000, //   ███   
		8'b01000100, //  █   █  
		8'b00000100, //      █
		8'b00111000, //   ███
		8'b00000100, //      █
		8'b01111100, //  ████
		8'b00000000, //
		
		8'b00000000, //
		8'b00001100, //     ██
		8'b00010100, //    █ █
		8'b00100100, //   █  █
		8'b01111100, //  █████
		8'b00000100, //      █
		8'b00000100, //      █
		8'b00000000, //
	
		8'b00000000, //
		8'b01111000, //  ████   
		8'b01000000, //  █
		8'b01110000, //  ███
		8'b00001000, //     █
		8'b01001000, //  █  █
		8'b01110000, //  ███
		8'b00000000, //
		
		8'b00000000, //
		8'b00111100, //   ████ 
		8'b01000000, //  █
		8'b01111000, //  ████ 
		8'b01000100, //  █   █
		8'b01000100, //  █   █
		8'b00111000, //   ███
		8'b00000000, //
		
		8'b00000000, //
		8'b01111110, //  ██████ 
		8'b00000010, //       █
		8'b00000100, //      █
		8'b00001000, //     █
		8'b00010000, //    █
		8'b00010000, //    █
		8'b00000000, //  

		8'b00000000, //
		8'b00111000, //   ███   
		8'b01000100, //  █   █ 
		8'b01000100, //  █   █
		8'b00111000, //   ███ 
		8'b01000100, //  █   █ 
		8'b01111100, //  █████ 
		8'b00000000, //
		
		8'b00000000, //
		8'b00110000, //   ██     
		8'b01001000, //  █  █   
		8'b01001000, //  █  █ 
		8'b00111000, //   ███  
		8'b00001000, //     █
		8'b00001000, //     █
		8'b00000000, //
		
	};
	
	assign data = ROM[address];

endmodule 